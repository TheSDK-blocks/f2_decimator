../../../TheSDK_generators/verilog/tb_f2_decimator.v