../../../TheSDK_generators/verilog/f2_decimator.v